module negate_32(A, S);
        
    input [31:0] A;

    output [31:0] S;

    not not_0(S[0], A[0]);
    not not_1(S[1], A[1]);
    not not_2(S[2], A[2]);
    not not_3(S[3], A[3]);
    not not_4(S[4], A[4]);
    not not_5(S[5], A[5]);
    not not_6(S[6], A[6]);
    not not_7(S[7], A[7]);
    not not_8(S[8], A[8]);
    not not_9(S[9], A[9]);
    not not_10(S[10], A[10]);
    not not_11(S[11], A[11]);
    not not_12(S[12], A[12]);
    not not_13(S[13], A[13]);
    not not_14(S[14], A[14]);
    not not_15(S[15], A[15]);
    not not_16(S[16], A[16]);
    not not_17(S[17], A[17]);
    not not_18(S[18], A[18]);
    not not_19(S[19], A[19]);
    not not_20(S[20], A[20]);
    not not_21(S[21], A[21]);
    not not_22(S[22], A[22]);
    not not_23(S[23], A[23]);
    not not_24(S[24], A[24]);
    not not_25(S[25], A[25]);
    not not_26(S[26], A[26]);
    not not_27(S[27], A[27]);
    not not_28(S[28], A[28]);
    not not_29(S[29], A[29]);
    not not_30(S[30], A[30]);
    not not_31(S[31], A[31]);

endmodule